// This file sets values for constants that may be affected by parameter values
  parameter [15:0] SAMPLE_SIZE  = 16'h0200;
  parameter [15:0] SAMPLING_FREQUENCY  = 16'h0400;
  parameter [15:0] NUM_TRAIN_CELLS  = 16'h000c;
  parameter [15:0] NUM_GUARD_CELLS  = 16'h0004;
  parameter [15:0] THRESHOLD_FACTOR  = 16'h0005;
  parameter [0:0] ocpi_debug  = 1'b0;
  parameter [1:0] ocpi_endian  = 2'b00;
  parameter [7:0] ocpi_version  = 8'h02;
  parameter [7:0] ocpi_max_opcode_input  = 8'h00;
  parameter [31:0] ocpi_max_bytes_input  = 32'h00002000;
  parameter [7:0] ocpi_max_opcode_output  = 8'h00;
  parameter [31:0] ocpi_max_bytes_output  = 32'h00002000;
  parameter [15:0] ocpi_max_latency_output  = 16'h0100;
  localparam ocpi_buffer_size_output_offset = 0;
  localparam ocpi_buffer_size_output_nbytes_1 = 1;
  localparam ocpi_blocked_output_offset = 4;
  localparam ocpi_blocked_output_nbytes_1 = 3;
  localparam ocpi_latency_output_offset = 8;
  localparam ocpi_latency_output_nbytes_1 = 1;
  localparam ocpi_messages_output_offset = 12;
  localparam ocpi_messages_output_nbytes_1 = 3;
  localparam ocpi_bytes_output_offset = 16;
  localparam ocpi_bytes_output_nbytes_1 = 3;
  localparam ocpi_sizeof_non_raw_properties = 20;
localparam ocpi_port_ctl_MAddr_width = 5;
localparam ocpi_port_ctl_MData_width = 32;
localparam ocpi_port_ctl_MByteEn_width = 4;
localparam ocpi_port_input_MData_width = 32;
localparam ocpi_port_input_MByteEn_width = 1;
localparam ocpi_port_input_MDataInfo_width = 1;
localparam ocpi_port_input_data_width = 32;
localparam ocpi_port_input_byte_width = 32;
localparam ocpi_port_output_MData_width = 32;
localparam ocpi_port_output_MByteEn_width = 1;
localparam ocpi_port_output_MDataInfo_width = 1;
localparam ocpi_port_output_data_width = 32;
localparam ocpi_port_output_byte_width = 32;

